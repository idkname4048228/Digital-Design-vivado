`timescale 1ns / 10ps
module Top();
    reg  A[3:0];
    wire B[7:0];
    wire C[7:0];

    
    initial begin
        #50
            A[0] = 1'b0;
            A[1] = 1'b0;
            A[2] = 1'b0;
            A[3] = 1'b0;
        #50
            A[0] = 1'b1;
        #50
            A[0] = 1'b0;
            A[1] = 1'b1;
        #50
            A[0] = 1'b1;
        #50
            A[0] = 1'b0;
            A[1] = 1'b0;
            A[2] = 1'b1;
        #50
            A[0] = 1'b1;
        #50
            A[0] = 1'b0;
            A[1] = 1'b1;
        #50
            A[0] = 1'b1;
        
        #50
            A[0] = 1'b0;
            A[1] = 1'b0;
            A[2] = 1'b0;
            A[3] = 1'b1;
        #50
            A[0] = 1'b1;
        #50
            A[0] = 1'b0;
            A[1] = 1'b1;
        #50
            A[0] = 1'b1;
        #50
            A[0] = 1'b0;
            A[1] = 1'b0;
            A[2] = 1'b1;
        #50
            A[0] = 1'b1;
        #50
            A[0] = 1'b0;
            A[1] = 1'b1;
        #50
            A[0] = 1'b1;
        #50 $finish;
    end
	

	four_to_sixteen_decoder u1(
        .A({A[3], A[2], A[1], A[0]}),//x, y, z
        .B({B[0], B[1], B[2], B[3], B[4], B[5], B[6], B[7]}),
        .C({C[0], C[1], C[2], C[3], C[4], C[5], C[6], C[7]})
    );

endmodule